library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.PACKAGE_MIPS.all;



ENTITY ADD4 IS 
 GENERIC(
         n:INTEGER
         );
 PORT(
		Xin		:IN		STD_LOGIC_VECTOR(n-1 DOWNTO 0):=(OTHERS=>'0');
		Sout	:OUT	STD_LOGIC_VECTOR(n-1 DOWNTO 0):=(OTHERS=>'0');
		Cout	:OUT	STD_LOGIC:='0'
      );
END ADD4;

ARCHITECTURE STRUCTURAL OF ADD4 IS 
  SIGNAL THREE 	:STD_LOGIC_VECTOR(n-1 DOWNTO 0);
  SIGNAL VDD	:STD_LOGIC:='1';
  SIGNAL GND	:STD_LOGIC:='0';
  SIGNAL CC		:STD_LOGIC_VECTOR(n-1 DOWNTO 2):=(OTHERS=>'0');
 BEGIN
 THREE<=CC&VDD&VDD;
 
G:CPA_FA GENERIC MAP (n) PORT MAP (Xin,THREE,VDD,Sout,Cout);


END STRUCTURAL;
