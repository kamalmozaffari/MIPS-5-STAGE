library ieee;
use ieee.std_logic_1164.all;
USE WORK.PACKAGE_MIPS.ALL;

ENTITY ALU IS
GENERIC (
		n:integer
	);
PORT(
	INPUT_1		:IN		STD_LOGIC_VECTOR(n-1	DOWNTO 0):=(OTHERS=>'0');
    INPUT_2		:IN		STD_LOGIC_VECTOR(n-1 	DOWNTO 0):=(OTHERS=>'0');
    AluOp		:IN		STD_LOGIC_VECTOR(1		DOWNTO 0):=(OTHERS=>'0');
	DATA_OUT	:OUT	STD_LOGIC_VECTOR(n-1	DOWNTO 0):=(OTHERS=>'0');
	carry		:OUT	STD_LOGIC
		);
end;

Architecture ST of ALU is 
SIGNAL R_AND_S,R_XOR_S,NOT_INPUT_2,IN_ADD_SUB,ADD_SUB	:STD_LOGIC_VECTOR(n-1 DOWNTO 0):=(OTHERS=>'0');
begin --architecture
NOT_INPUT_2	<= NOT(INPUT_2);
R_AND_S		<=INPUT_1 AND INPUT_2;
R_XOR_S		<=INPUT_1 XOR INPUT_2;

G_MUX2TO1		:	MUX2TO1		GENERIC MAP(n)		PORT MAP	(INPUT_2,NOT_INPUT_2,AluOp(0),IN_ADD_SUB);
G_ADDER_SUBTRUCT:	CPA_FA	GENERIC MAP	(n) PORT MAP 	(INPUT_1,IN_ADD_SUB,AluOp(0),ADD_SUB,carry);
G_MUX4TO1		:	MUX4TO1 GENERIC MAP (n) PORT MAP 	(ADD_SUB,ADD_SUB,R_AND_S,R_XOR_S,AluOp,DATA_OUT);



END ARCHITECTURE;